

module Top
   ()

endmodule