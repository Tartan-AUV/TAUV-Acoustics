

module top_pl
   (output reg AFE0_DIR);

endmodule
